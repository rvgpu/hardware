`define OPCODE_ADD 8'h01
`define OPCODE_SUB 8'h02